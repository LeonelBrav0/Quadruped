module tb_ne_write_coeff_buffer();

endmodule