interface kria_kr260_IO;
    logic 

endinterface