//--------------------------------------------------------------------------
//
//          PROJECT N: AXI4_LITE NEURAL ENGINE
//
//--------------------------------------------------------------------------
//
//  File: hw_ne_arbiter.sv
//  
//  Author: Marc Francis Leonel Bravo
//
//--------------------------------------------------------------------------
//
//  Abstract    :   Hardware arbitration for coeff buffer spsram banks
//
//--------------------------------------------------------------------------
//  Revision History
//  @ 09/29/2023    :   initial
//  Initial commit
//--------------------------------------------------------------------------