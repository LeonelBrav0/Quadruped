module q_top_tb();


reg  [15:0] a;
reg  [15:0] b;
wire [15:0] c;

initial begin
    $display("HELLO WORLD TESTBENCH");
end



endmodule