module q_top(
    p_fan_en_b,
    p_pmod1,
    p_pmod2,
    p_pmod3,
    p_pmod4,
    p_rpi_header
);



endmodule

